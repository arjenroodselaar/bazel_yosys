version https://git-lfs.github.com/spec/v1
oid sha256:739edd0f0b073a723f058b89c917fd59b642443224094989af603cd621e52c72
size 30744
