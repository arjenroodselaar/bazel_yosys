version https://git-lfs.github.com/spec/v1
oid sha256:cfc8756b1cd925a8dfa7b395ed086558768a926dd44e72d5490f6db0b9bf6883
size 39800
