version https://git-lfs.github.com/spec/v1
oid sha256:f93778126355215298683d50035f61de9958f4efc0ed0bab51d4559b913a1a5d
size 50688
