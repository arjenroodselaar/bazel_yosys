version https://git-lfs.github.com/spec/v1
oid sha256:8b0b0c821b4ea6e40e5e8b38d2f88caed42453c9eb259cd31a0c8844d862020f
size 4096
