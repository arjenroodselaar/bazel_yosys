version https://git-lfs.github.com/spec/v1
oid sha256:1ef3c5fda008b7412d9b8c53b641d76509b22236b191dbbae255f0565f60cf2d
size 2048
