version https://git-lfs.github.com/spec/v1
oid sha256:3029063c475a211f980a0eb590cdb4dfa2d6055bdb2c2ab4956017efe248579e
size 812
