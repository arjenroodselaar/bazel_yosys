version https://git-lfs.github.com/spec/v1
oid sha256:b9237fb2badbc9e1640c1d2e98591f1d19e066cb2caee3a406de84a8445e5ed0
size 1801
