`define RISCV_FORMAL
`define RISCV_FORMAL_NRET 1
`define RISCV_FORMAL_XLEN 32
`define RISCV_FORMAL_ILEN 32
`define RISCV_FORMAL_RESET_CYCLES 1
`define RISCV_FORMAL_CHECK_CYCLE 20
`define RISCV_FORMAL_CHANNEL_IDX 0
`define RISCV_FORMAL_CSR_MCYCLE
`define RISCV_FORMAL_CSR_MINSTRET
`define RISCV_FORMAL_COMPRESSED
`define RISCV_FORMAL_ALIGNED_MEM
`define RISCV_FORMAL_ALTOPS
`define PICORV32_CSR_RESTRICT
`define PICORV32_TESTBUG_NONE
`define DEBUGNETS
`include "hdl/cpu/riscv_formal/checks/rvfi_macros.vh"
