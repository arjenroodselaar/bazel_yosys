version https://git-lfs.github.com/spec/v1
oid sha256:184031b7cc919da2200909731491cae24cda67283738bcd5b5edf435381674b4
size 846
