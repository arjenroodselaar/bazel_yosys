version https://git-lfs.github.com/spec/v1
oid sha256:c0837dc7752f55d523de75f204b973118061f990cef6db89ccf3ef387460754d
size 1024
