version https://git-lfs.github.com/spec/v1
oid sha256:26ba71d1655fe69195e4f4fa6200e3330c250fdc4453c57036f727a298743b47
size 165200
