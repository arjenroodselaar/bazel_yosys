version https://git-lfs.github.com/spec/v1
oid sha256:e5a598328ab3d53ffe49f362ed559cce3de97347f7b7be1cd45a20d7daadde25
size 6129
