version https://git-lfs.github.com/spec/v1
oid sha256:52b6b32e947e0d3c986e4373dd5bc5fd5cad3a31598629238f7741242c50ef87
size 81600
