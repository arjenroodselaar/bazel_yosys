version https://git-lfs.github.com/spec/v1
oid sha256:3806f41b17faadfe54a717655347690e91d2232f74509ee937ddd0d255490133
size 939
