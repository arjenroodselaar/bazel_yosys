version https://git-lfs.github.com/spec/v1
oid sha256:8fe7addb93b1effe33b19dacbbeca754b18d224de786769a7b7a99464f407e68
size 50688
