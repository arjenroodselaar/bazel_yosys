version https://git-lfs.github.com/spec/v1
oid sha256:279b32864ddc83716a70c0fb055ecb1d5947b8bf0903f547d9fb48fb95f25405
size 50688
