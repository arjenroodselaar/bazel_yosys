version https://git-lfs.github.com/spec/v1
oid sha256:d04a280346b303e0ae90b0abfd936828d28dce3fd103848a0b77fe58d1344dde
size 949
