version https://git-lfs.github.com/spec/v1
oid sha256:b56c162108bbaff9887cb7cf788444b295388402bc5b707c570007123fe34748
size 1748
