version https://git-lfs.github.com/spec/v1
oid sha256:71964f2aab79035acd9813f18b7c747e678eedaf1bdd28755df02c7e135eef6f
size 801
