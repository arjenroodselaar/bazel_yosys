version https://git-lfs.github.com/spec/v1
oid sha256:a1e5162547680cec95ead184583f3f00d8410417d6a308b95e2eb218efb7a74b
size 900
