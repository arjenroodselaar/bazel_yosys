version https://git-lfs.github.com/spec/v1
oid sha256:759306a7e7df71609beacae9fae2a423192c84b7bca4e4fcc8d325ece8a73d7d
size 1174
