version https://git-lfs.github.com/spec/v1
oid sha256:14c8c92057d492b9aa009c802347a3b0bf5d38ddf20e487f482713b8e1de9251
size 59136
